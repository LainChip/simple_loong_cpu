// TODO: XRB