module scoreboard(
    input reg_0,
    input reg_1,
    input reg_2,
    input reg_3,


);

endmodule