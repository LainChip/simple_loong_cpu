`ifndef _TLB_HEADER
`define _TLB_HEADER

/*--JSON--{"module_name":"deperated","module_ver":"3","module_type":"module"}--JSON--*/
`endif
