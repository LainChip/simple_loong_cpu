`include "common.svh"
`include "decoder.svh"
`include "tlb.svh"

`ifdef _TLB_VER_1

module tlb(

);

endmodule : tlb

`endif 