/*
2023-1 v1
*/

module divider (
    input clk,
    input rst_n,

    input  div_signed_i,
    input  [31:0] Z_i,
    input  [31:0] D_i,
    output [31:0] q_o, s_o
);



endmodule