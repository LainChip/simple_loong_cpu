`include "decoder.svh"
/*--JSON--{"module_name":"scoreboard","module_ver":"2","module_type":"module"}--JSON--*/
module issue(
    input logic clk,
    input logic rst_n,
    input inst_t[1:0] inst,

);
endmodule