`include "common.svh"
`include "lsu_types.svh"

module lsu_test_plantform (
	input clk,    // Clock
	input rst_n  // Asynchronous reset active low
;

endmodule : lsu_test_plantform