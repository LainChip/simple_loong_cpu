`ifndef _COMMON_HEADER
`define _COMMON_HEADER

`timescale 1ns/1ps

`define __AXI_CONVERTER_VER_1

`define _CACHE_BUS_DATA_LEN (32)

`endif
