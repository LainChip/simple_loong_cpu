`include "common.svh"
`include "decoder.svh"

module decoder(
    input logic[31:0] inst_i,
    output decode_info_t decode_info_o,
    output logic[31:0][7:0] inst_string_o
);

    always_comb begin
        casez(inst_i)
            32'b010011??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = `_BRANCH_INDIRECT;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_BPF;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = `_USE_EX;
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd106 ,8'd105 ,8'd114 ,8'd108}; //jirl
            end
            32'b010100??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = `_BRANCH_IMMEDIATE;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                inst_string_o = {8'd98}; //b
            end
            32'b010101??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = `_BRANCH_IMMEDIATE;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd1;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_BPF;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_BL;
                inst_string_o = {8'd98 ,8'd108}; //bl
            end
            32'b010110??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_EQL;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                inst_string_o = {8'd98 ,8'd101 ,8'd113}; //beq
            end
            32'b010111??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_NEQ;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                inst_string_o = {8'd98 ,8'd110 ,8'd101}; //bne
            end
            32'b011000??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_LSS;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                inst_string_o = {8'd98 ,8'd108 ,8'd116}; //blt
            end
            32'b011001??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_GER;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                inst_string_o = {8'd98 ,8'd103 ,8'd101}; //bge
            end
            32'b011010??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_LTU;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                inst_string_o = {8'd98 ,8'd108 ,8'd116 ,8'd117}; //bltu
            end
            32'b011011??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_GEU;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                inst_string_o = {8'd98 ,8'd103 ,8'd101 ,8'd117}; //bgeu
            end
            32'b0001010?????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_LUI;
                decode_info_o.ex.opd_type = `_OPD_IMM_S20;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_W;
                inst_string_o = {8'd108 ,8'd117 ,8'd49 ,8'd50 ,8'd105 ,8'd46 ,8'd119}; //lu12i.w
            end
            32'b0001110?????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_ADD;
                decode_info_o.ex.opd_type = `_OPD_IMM_S20;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_W;
                inst_string_o = {8'd112 ,8'd99 ,8'd97 ,8'd100 ,8'd100 ,8'd117 ,8'd49 ,8'd50 ,8'd105}; //pcaddu12i
            end
            32'b00000100????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd1;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_CSR;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_M2,`_USE_M2};
                decode_info_o.is.reg_type = `_REG_TYPE_CSRXCHG;
                inst_string_o = {8'd99 ,8'd115 ,8'd114 ,8'd119 ,8'd114 ,8'd120 ,8'd99 ,8'd104 ,8'd103}; //csrwrxchg
            end
            32'b0000001000??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info_o.ex.opd_type = `_OPD_IMM_S12;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd115 ,8'd108 ,8'd116 ,8'd105}; //slti
            end
            32'b0000001001??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info_o.ex.opd_type = `_OPD_IMM_S12;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd115 ,8'd108 ,8'd116 ,8'd117 ,8'd105}; //sltui
            end
            32'b0000001010??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_ADD;
                decode_info_o.ex.opd_type = `_OPD_IMM_S12;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd97 ,8'd100 ,8'd100 ,8'd105 ,8'd46 ,8'd119}; //addi.w
            end
            32'b0000001101??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_AND;
                decode_info_o.ex.opd_type = `_OPD_IMM_U12;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd97 ,8'd110 ,8'd100 ,8'd105}; //andi
            end
            32'b0000001110??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_OR;
                decode_info_o.ex.opd_type = `_OPD_IMM_U12;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd111 ,8'd114 ,8'd105}; //ori
            end
            32'b0000001111??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_XOR;
                decode_info_o.ex.opd_type = `_OPD_IMM_U12;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd120 ,8'd111 ,8'd114 ,8'd105}; //xori
            end
            32'b0010100000??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_BYTE;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd108 ,8'd100 ,8'd46 ,8'd98}; //ld.b
            end
            32'b0010100001??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_HALF;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd108 ,8'd100 ,8'd46 ,8'd104}; //ld.h
            end
            32'b0010100010??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd108 ,8'd100 ,8'd46 ,8'd119}; //ld.w
            end
            32'b0010100100??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_BYTE;
                decode_info_o.m1.mem_write = 1'd1;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                inst_string_o = {8'd115 ,8'd116 ,8'd46 ,8'd98}; //st.b
            end
            32'b0010100101??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_HALF;
                decode_info_o.m1.mem_write = 1'd1;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                inst_string_o = {8'd115 ,8'd116 ,8'd46 ,8'd104}; //st.h
            end
            32'b0010100110??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info_o.m1.mem_write = 1'd1;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                inst_string_o = {8'd115 ,8'd116 ,8'd46 ,8'd119}; //st.w
            end
            32'b0010101000??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_UBYTE;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd108 ,8'd100 ,8'd46 ,8'd98 ,8'd117}; //ld.bu
            end
            32'b0010101001??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_UHALF;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd108 ,8'd100 ,8'd46 ,8'd104 ,8'd117}; //ld.hu
            end
            32'b0010101010??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_UWORD;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd108 ,8'd100 ,8'd46 ,8'd119 ,8'd117}; //ld.wu
            end
            32'b00000000000100000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_ADD;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd97 ,8'd100 ,8'd100 ,8'd46 ,8'd119}; //add.w
            end
            32'b00000000000100010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_SUB;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd115 ,8'd117 ,8'd98 ,8'd46 ,8'd119}; //sub.w
            end
            32'b00000000000100100???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd115 ,8'd108 ,8'd116}; //slt
            end
            32'b00000000000100101???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd115 ,8'd108 ,8'd116 ,8'd117}; //sltu
            end
            32'b00000000000101000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_NOR;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd110 ,8'd111 ,8'd114}; //nor
            end
            32'b00000000000101001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_AND;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd97 ,8'd110 ,8'd100}; //and
            end
            32'b00000000000101010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_OR;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd111 ,8'd114}; //or
            end
            32'b00000000000101011???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_XOR;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd120 ,8'd111 ,8'd114}; //xor
            end
            32'b00000000000101110???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_SL;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd115 ,8'd108 ,8'd108 ,8'd46 ,8'd119}; //sll.w
            end
            32'b00000000000101111???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_SR;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd115 ,8'd114 ,8'd108 ,8'd46 ,8'd119}; //srl.w
            end
            32'b00000000000110000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_SR;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd115 ,8'd114 ,8'd97 ,8'd46 ,8'd119}; //sra.w
            end
            32'b00000000000111000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_MUL;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd109 ,8'd117 ,8'd108 ,8'd46 ,8'd119}; //mul.w
            end
            32'b00000000000111001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_MULH;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd109 ,8'd117 ,8'd108 ,8'd104 ,8'd46 ,8'd119}; //mulh.w
            end
            32'b00000000000111010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_MULH;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd109 ,8'd117 ,8'd108 ,8'd104 ,8'd46 ,8'd119 ,8'd117}; //mulh.wu
            end
            32'b00000000001000000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_DIV;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd100 ,8'd105 ,8'd118 ,8'd46 ,8'd119}; //div.w
            end
            32'b00000000001000001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_MOD;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd109 ,8'd111 ,8'd100 ,8'd46 ,8'd119}; //mod.w
            end
            32'b00000000001000010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_DIV;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd100 ,8'd105 ,8'd118 ,8'd46 ,8'd119 ,8'd117}; //div.wu
            end
            32'b00000000001000011???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_MOD;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                inst_string_o = {8'd109 ,8'd111 ,8'd100 ,8'd46 ,8'd119 ,8'd117}; //mod.wu
            end
            32'b00000000001010100???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_SYSCALL;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                inst_string_o = {8'd98 ,8'd114 ,8'd101 ,8'd97 ,8'd107}; //break
            end
            32'b00000000001010110???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_SYSCALL;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                inst_string_o = {8'd115 ,8'd121 ,8'd115 ,8'd99 ,8'd97 ,8'd108 ,8'd108}; //syscall
            end
            32'b00000000010000001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_SL;
                decode_info_o.ex.opd_type = `_OPD_IMM_U5;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd115 ,8'd108 ,8'd108 ,8'd105 ,8'd46 ,8'd119}; //slli.w
            end
            32'b00000000010001001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_SR;
                decode_info_o.ex.opd_type = `_OPD_IMM_U5;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd115 ,8'd114 ,8'd108 ,8'd105 ,8'd46 ,8'd119}; //srli.w
            end
            32'b00000000010010001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = `_ALU_TYPE_SR;
                decode_info_o.ex.opd_type = `_OPD_IMM_U5;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b0;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd115 ,8'd114 ,8'd97 ,8'd105 ,8'd46 ,8'd119}; //srai.w
            end
            32'b00000110010010001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                inst_string_o = {8'd105 ,8'd100 ,8'd108 ,8'd101}; //idle
            end
            32'b00000110010010011???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd1;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_M2,`_USE_M2};
                decode_info_o.is.reg_type = `_REG_TYPE_INVTLB;
                inst_string_o = {8'd105 ,8'd110 ,8'd118 ,8'd116 ,8'd108 ,8'd98}; //invtlb
            end
            32'b0000000000000000011000??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd1;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_CSR;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RDCNTID;
                inst_string_o = {8'd114 ,8'd100 ,8'd99 ,8'd110 ,8'd116 ,8'd105 ,8'd100 ,8'd46 ,8'd119}; //rdcntid.w
            end
            32'b0000000000000000011000??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_LOW;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_CSR;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd114 ,8'd100 ,8'd99 ,8'd110 ,8'd116 ,8'd118 ,8'd108 ,8'd46 ,8'd119}; //rdcntvl.w
            end
            32'b0000000000000000011001??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_HIGH;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_CSR;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd114 ,8'd100 ,8'd99 ,8'd110 ,8'd116 ,8'd118 ,8'd104 ,8'd46 ,8'd119}; //rdcntvh.w
            end
            32'b0000011001001000001010??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd1;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd116 ,8'd108 ,8'd98 ,8'd115 ,8'd114 ,8'd99 ,8'd104}; //tlbsrch
            end
            32'b0000011001001000001011??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd1;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd116 ,8'd108 ,8'd98 ,8'd114 ,8'd100}; //tlbrd
            end
            32'b0000011001001000001100??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd1;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd116 ,8'd108 ,8'd98 ,8'd119 ,8'd114}; //tlbwr
            end
            32'b0000011001001000001101??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd1;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                inst_string_o = {8'd116 ,8'd108 ,8'd98 ,8'd102 ,8'd105 ,8'd108 ,8'd108}; //tlbfill
            end
            32'b0000011001001000001110??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd1;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                inst_string_o = {8'd101 ,8'd114 ,8'd116 ,8'd110}; //ertn
            end
            default: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m2.rdcntv_type = `_RDCNTV_TYPE_NONE;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_INVALID;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m1.tlbwr_en = 1'd0;
                decode_info_o.m1.tlbfill_en = 1'd0;
                decode_info_o.m1.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = 4'b1111;
                inst_string_o = {8'd78 ,8'd79 ,8'd78 ,8'd69 ,8'd86 ,8'd65 ,8'd76 ,8'd73 ,8'd68}; //NONEVALID
            end
        endcase
    end

endmodule
