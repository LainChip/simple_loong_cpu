`ifndef _TLB_HEADER
`define _TLB_HEADER

`endif
