`ifndef _BPU_SVH_
`define _BPU_SVH_

`define SCS_STRONGLY_TAKEN 2'b11
`define SCS_WEAKLY_TAKEN 2'b10
`define SCS_WEAKLY_NOT_TAKEN 2'b01
`define SCS_STRONGLY_NOT_TAKEN 2'b00

`define SCS_STRONGLY_GLOBAL 2'b11
`define SCS_WEAKLY_GLOBAL 2'b10
`define SCS_WEAKLY_LOCAL 2'b01
`define SCS_STRONGLY_LOCAL 2'b00

























`endif // _BPU_SVH_