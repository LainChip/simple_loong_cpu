`include "common.svh"
`include "decoder.svh"

module decoder(
    input logic[31:0] inst_i,
    input logic fetch_err_i,
    output decode_info_t decode_info_o,
    output logic[31:0][7:0] inst_string_o
);

    always_comb begin
        unique casez(inst_i)
            32'b010011??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = `_BRANCH_INDIRECT;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S16;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_LI;
                decode_info_o.m2.alu_op = `_ALU_STYPE_PCPLUS4;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //jirl
            end
            32'b010100??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = `_BRANCH_INDIRECT;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S26;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //b
            end
            32'b010101??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = `_BRANCH_INDIRECT;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_BL1;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S26;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_LI;
                decode_info_o.m2.alu_op = `_ALU_STYPE_PCPLUS4;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //bl
            end
            32'b010110??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = `_BRANCH_CONDITION;
                decode_info_o.m1.cmp_type = `_CMP_E;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RD;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S16;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //beq
            end
            32'b010111??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = `_BRANCH_CONDITION;
                decode_info_o.m1.cmp_type = `_CMP_NE;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RD;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S16;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //bne
            end
            32'b011000??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = `_BRANCH_CONDITION;
                decode_info_o.m1.cmp_type = `_CMP_LT;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RD;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S16;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //blt
            end
            32'b011001??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = `_BRANCH_CONDITION;
                decode_info_o.m1.cmp_type = `_CMP_GE;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RD;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S16;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //bge
            end
            32'b011010??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = `_BRANCH_CONDITION;
                decode_info_o.m1.cmp_type = `_CMP_LTU;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RD;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S16;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //bltu
            end
            32'b011011??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = `_BRANCH_CONDITION;
                decode_info_o.m1.cmp_type = `_CMP_GEU;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RD;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S16;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //bgeu
            end
            32'b0001010?????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_IMM;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_S20;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_LI;
                decode_info_o.m2.alu_op = `_ALU_STYPE_LUI;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //lu12i.w
            end
            32'b0001110?????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_IMM;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_S20;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_LI;
                decode_info_o.m2.alu_op = `_ALU_STYPE_PCADDUI;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //pcaddu12i
            end
            32'b00000100????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_CSR;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RD;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd1;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd1;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //csrwrxchg
            end
            32'b00100000????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd1;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd1;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S14;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //ll.w
            end
            32'b00100001????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info_o.m1.mem_write = 1'd1;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd1;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RD;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S14;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //sc.w
            end
            32'b0000001000??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_IMM;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_S12;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_CMP;
                decode_info_o.m2.alu_op = `_ALU_STYPE_SLT;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //slti
            end
            32'b0000001001??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_IMM;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_S12;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_CMP;
                decode_info_o.m2.alu_op = `_ALU_STYPE_SLTU;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //sltui
            end
            32'b0000001010??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_IMM;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_S12;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_INT;
                decode_info_o.m2.alu_op = `_ALU_STYPE_ADD;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //addi.w
            end
            32'b0000001101??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_IMM;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U12;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_BW;
                decode_info_o.m2.alu_op = `_ALU_STYPE_AND;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //andi
            end
            32'b0000001110??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_IMM;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U12;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_BW;
                decode_info_o.m2.alu_op = `_ALU_STYPE_OR;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //ori
            end
            32'b0000001111??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_IMM;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U12;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_BW;
                decode_info_o.m2.alu_op = `_ALU_STYPE_XOR;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //xori
            end
            32'b0000011000??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = `_MEM_TYPE_BYTE;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd1;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd1;
                decode_info_o.m1.refetch = 1'd1;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //cacop
            end
            32'b0010100000??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = `_MEM_TYPE_BYTE;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd1;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //ld.b
            end
            32'b0010100001??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = `_MEM_TYPE_HALF;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd1;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //ld.h
            end
            32'b0010100010??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd1;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //ld.w
            end
            32'b0010100100??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = `_MEM_TYPE_BYTE;
                decode_info_o.m1.mem_write = 1'd1;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RD;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //st.b
            end
            32'b0010100101??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = `_MEM_TYPE_HALF;
                decode_info_o.m1.mem_write = 1'd1;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RD;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //st.h
            end
            32'b0010100110??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info_o.m1.mem_write = 1'd1;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RD;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //st.w
            end
            32'b0010101000??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = `_MEM_TYPE_UBYTE;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd1;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //ld.bu
            end
            32'b0010101001??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = `_MEM_TYPE_UHALF;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd1;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_ADDR_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //ld.hu
            end
            32'b0010101011??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //preld_nop
            end
            32'b00000000000100000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_INT;
                decode_info_o.m2.alu_op = `_ALU_STYPE_ADD;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //add.w
            end
            32'b00000000000100010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_INT;
                decode_info_o.m2.alu_op = `_ALU_STYPE_SUB;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //sub.w
            end
            32'b00000000000100100???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_CMP;
                decode_info_o.m2.alu_op = `_ALU_STYPE_SLT;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //slt
            end
            32'b00000000000100101???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'd1;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'd1;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_CMP;
                decode_info_o.m2.alu_op = `_ALU_STYPE_SLTU;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //sltu
            end
            32'b00000000000101000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_BW;
                decode_info_o.m2.alu_op = `_ALU_STYPE_NOR;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //nor
            end
            32'b00000000000101001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_BW;
                decode_info_o.m2.alu_op = `_ALU_STYPE_AND;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //and
            end
            32'b00000000000101010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_BW;
                decode_info_o.m2.alu_op = `_ALU_STYPE_OR;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //or
            end
            32'b00000000000101011???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = `_FUSEL_EX_ALU;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_BW;
                decode_info_o.m2.alu_op = `_ALU_STYPE_XOR;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //xor
            end
            32'b00000000000101110???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_SFT;
                decode_info_o.m2.alu_op = `_ALU_STYPE_SLL;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //sll.w
            end
            32'b00000000000101111???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_SFT;
                decode_info_o.m2.alu_op = `_ALU_STYPE_SRL;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //srl.w
            end
            32'b00000000000110000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_SFT;
                decode_info_o.m2.alu_op = `_ALU_STYPE_SRA;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //sra.w
            end
            32'b00000000000111000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'd1;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_MUL;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = `_MUL_TYPE_MULL;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //mul.w
            end
            32'b00000000000111001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'd1;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_MUL;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = `_MUL_TYPE_MULH;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //mulh.w
            end
            32'b00000000000111010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'd1;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_MUL;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = `_MUL_TYPE_MULHU;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //mulh.wu
            end
            32'b00000000001000000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'd1;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = `_FUSEL_WB_DIV;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = `_DIV_TYPE_DIV;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //div.w
            end
            32'b00000000001000001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'd1;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = `_FUSEL_WB_DIV;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = `_DIV_TYPE_MOD;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //mod.w
            end
            32'b00000000001000010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'd1;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = `_FUSEL_WB_DIV;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = `_DIV_TYPE_DIVU;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //div.wu
            end
            32'b00000000001000011???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'd1;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'd1;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'd1;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = `_FUSEL_WB_DIV;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = `_DIV_TYPE_MODU;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //mod.wu
            end
            32'b00000000001010110???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd1;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //syscall
            end
            32'b00000000001010110???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd1;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //break
            end
            32'b00000000010000001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_IMM;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_SFT;
                decode_info_o.m2.alu_op = `_ALU_STYPE_SLL;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //slli.w
            end
            32'b00000000010001001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_IMM;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_SFT;
                decode_info_o.m2.alu_op = `_ALU_STYPE_SRL;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //srli.w
            end
            32'b00000000010010001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = `_FUSEL_M1_ALU;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_ALU;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_IMM;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = `_ALU_GTYPE_SFT;
                decode_info_o.m2.alu_op = `_ALU_STYPE_SRA;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //srai.w
            end
            32'b00000110010010001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd1;
                decode_info_o.m1.refetch = 1'd1;
                decode_info_o.m1.wait_inst = 1'd1;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //idle
            end
            32'b00000110010010011???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'd1;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_RK;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd1;
                decode_info_o.m1.refetch = 1'd1;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd1;
                inst_string_o = '0; //invtlb
            end
            32'b00111000011100100???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd1;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //dbar
            end
            32'b00111000011100101???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd1;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd1;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //ibar
            end
            32'b0000000000000000011000??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'd1;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_CSR;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_RJ;
                decode_info_o.is.reg_type_w = `_REG_W_RJD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //rdcnt.w
            end
            32'b0000000000000000011001??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = `_FUSEL_M2_CSR;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_RJD;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //rdcnth.w
            end
            32'b0000011001001000001010??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd1;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd1;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //tlbsrch
            end
            32'b0000011001001000001011??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd1;
                decode_info_o.m1.refetch = 1'd1;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd1;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //tlbrd
            end
            32'b0000011001001000001100??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd1;
                decode_info_o.m1.refetch = 1'd1;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd1;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //tlbwr
            end
            32'b0000011001001000001101??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd1;
                decode_info_o.m1.refetch = 1'd1;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd1;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //tlbfill
            end
            32'b0000011001001000001110??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.m2.need_csr = 1'b0;
                decode_info_o.m2.need_mul = 1'b0;
                decode_info_o.m2.need_div = 1'b0;
                decode_info_o.m2.need_lsu = 1'b0;
                decode_info_o.m2.need_bpu = 1'b0;
                decode_info_o.ex.latest_r0_ex = 1'b0;
                decode_info_o.m1.latest_r0_m1 = 1'b0;
                decode_info_o.m2.latest_r0_m2 = 1'b0;
                decode_info_o.wb.latest_r0_wb = 1'b0;
                decode_info_o.ex.latest_r1_ex = 1'b0;
                decode_info_o.m1.latest_r1_m1 = 1'b0;
                decode_info_o.m2.latest_r1_m2 = 1'b0;
                decode_info_o.wb.latest_r1_wb = 1'b0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = `_REG_R0_NONE;
                decode_info_o.is.reg_type_r1 = `_REG_R1_NONE;
                decode_info_o.is.reg_type_w = `_REG_W_NONE;
                decode_info_o.is.imm_type = `_IMM_U5;
                decode_info_o.ex.addr_imm_type = `_IMM_S12;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd1;
                decode_info_o.m1.priv_inst = 1'd1;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = '0; //ertn
            end
            default: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_read = 1'd0;
                decode_info_o.m2.mem_cacop = 1'd0;
                decode_info_o.m2.llsc_inst = 1'd0;
                decode_info_o.m1.ibarrier = 1'd0;
                decode_info_o.m1.dbarrier = 1'd0;
                decode_info_o.m1.branch_type = 2'd0;
                decode_info_o.m1.cmp_type = 3'd0;
                decode_info_o.wb.debug_inst = 32'd0;
                decode_info_o.m2.need_csr = 1'd0;
                decode_info_o.m2.need_mul = 1'd0;
                decode_info_o.m2.need_div = 1'd0;
                decode_info_o.m2.need_lsu = 1'd0;
                decode_info_o.m2.need_bpu = 1'd0;
                decode_info_o.ex.latest_r0_ex = 1'd0;
                decode_info_o.m1.latest_r0_m1 = 1'd0;
                decode_info_o.m2.latest_r0_m2 = 1'd0;
                decode_info_o.wb.latest_r0_wb = 1'd0;
                decode_info_o.ex.latest_r1_ex = 1'd0;
                decode_info_o.m1.latest_r1_m1 = 1'd0;
                decode_info_o.m2.latest_r1_m2 = 1'd0;
                decode_info_o.wb.latest_r1_wb = 1'd0;
                decode_info_o.ex.fu_sel_ex = 1'd0;
                decode_info_o.m1.fu_sel_m1 = 2'd0;
                decode_info_o.m2.fu_sel_m2 = 2'd0;
                decode_info_o.m2.fu_sel_wb = 1'd0;
                decode_info_o.is.reg_type_r0 = 2'd0;
                decode_info_o.is.reg_type_r1 = 1'd0;
                decode_info_o.is.reg_type_w = 2'd0;
                decode_info_o.is.imm_type = 3'd0;
                decode_info_o.ex.addr_imm_type = 2'd0;
                decode_info_o.m2.alu_grand_op = 2'd0;
                decode_info_o.m2.alu_op = 2'd0;
                decode_info_o.m1.ertn_inst = 1'd0;
                decode_info_o.m1.priv_inst = 1'd0;
                decode_info_o.m1.refetch = 1'd0;
                decode_info_o.m1.wait_inst = 1'd0;
                decode_info_o.m1.invalid_inst = 1'd0;
                decode_info_o.m1.syscall_inst = 1'd0;
                decode_info_o.m1.break_inst = 1'd0;
                decode_info_o.m2.csr_op_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                inst_string_o = {8'd78 ,8'd79 ,8'd78 ,8'd69 ,8'd86 ,8'd65 ,8'd76 ,8'd73 ,8'd68}; //NONEVALID
            end
        endcase
    end

endmodule
