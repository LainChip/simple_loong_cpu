/*
2023-1-17 v1
*/

// count leadding zero
