`include "common.svh"
`include "lsu_types.svh"

`ifdef __DLSU_VER_1

`endif