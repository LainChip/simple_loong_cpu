`include "common.svh"
`include "decoder.svh"

module(
    input logic[31:0] inst,
    output decode_info_t decode_info,
    output logic[31:0][7:0] inst_string
);

    always_comb begin
        casex(inst)
            32'b010011xxxxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = `_BRANCH_INDIRECT;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_EX;
                decode_info.is.use_time = `_USE_EX;
                decode_info.is.reg_type = `_REG_TYPE_RW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd106 ,8'd105 ,8'd114 ,8'd108}; //jirl
            end
            32'b010100xxxxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = `_BRANCH_IMMEDIATE;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_I;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd98}; //b
            end
            32'b010101xxxxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = `_BRANCH_IMMEDIATE;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_EX;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_BL;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd98 ,8'd108}; //bl
            end
            32'b010110xxxxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = `_BRANCH_CONDITION;
                decode_info.ex.cmp_type = `_CMP_EQL;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd98 ,8'd101 ,8'd113}; //beq
            end
            32'b010111xxxxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = `_BRANCH_CONDITION;
                decode_info.ex.cmp_type = `_CMP_NEQ;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd98 ,8'd110 ,8'd101}; //bne
            end
            32'b011000xxxxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = `_BRANCH_CONDITION;
                decode_info.ex.cmp_type = `_CMP_LSS;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd98 ,8'd108 ,8'd116}; //blt
            end
            32'b011001xxxxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = `_BRANCH_CONDITION;
                decode_info.ex.cmp_type = _CMP_GER;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd98 ,8'd103 ,8'd101}; //bge
            end
            32'b011010xxxxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = `_BRANCH_CONDITION;
                decode_info.ex.cmp_type = `_CMP_LTU;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd98 ,8'd108 ,8'd116 ,8'd117}; //bltu
            end
            32'b011011xxxxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = `_BRANCH_CONDITION;
                decode_info.ex.cmp_type = `_CMP_GEU;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd98 ,8'd103 ,8'd101 ,8'd117}; //bgeu
            end
            32'b0001010xxxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_LUI;
                decode_info.ex.opd_type = `_OPD_IMM_S20;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd108 ,8'd117 ,8'd49 ,8'd50 ,8'd105 ,8'd46 ,8'd119}; //lu12i.w
            end
            32'b0001110xxxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_ADD;
                decode_info.ex.opd_type = `_OPD_IMM_S20;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd112 ,8'd99 ,8'd97 ,8'd100 ,8'd100 ,8'd117 ,8'd49 ,8'd50 ,8'd105}; //pcaddu12i
            end
            32'b00000100xxxxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd1;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_M2,`_USE_M2};
                decode_info.is.reg_type = `_REG_TYPE_CSRXCHG;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd99 ,8'd115 ,8'd114 ,8'd120 ,8'd99 ,8'd104 ,8'd103}; //csrxchg
            end
            32'b0000001000xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info.ex.opd_type = `_OPD_IMM_S12;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd108 ,8'd116 ,8'd105}; //slti
            end
            32'b0000001001xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info.ex.opd_type = `_OPD_IMM_S12;
                decode_info.ex.opd_unsigned = 1'd1;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd108 ,8'd116 ,8'd117 ,8'd105}; //sltui
            end
            32'b0000001010xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_ADD;
                decode_info.ex.opd_type = `_OPD_IMM_S12;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd97 ,8'd100 ,8'd100 ,8'd105 ,8'd46 ,8'd119}; //addi.w
            end
            32'b0000001101xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_AND;
                decode_info.ex.opd_type = `_OPD_IMM_U12;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd97 ,8'd110 ,8'd100 ,8'd105}; //andi
            end
            32'b0000001110xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_OR;
                decode_info.ex.opd_type = `_OPD_IMM_U12;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd111 ,8'd114 ,8'd105}; //ori
            end
            32'b0000001111xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_XOR;
                decode_info.ex.opd_type = `_OPD_IMM_U12;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd120 ,8'd111 ,8'd114 ,8'd105}; //xori
            end
            32'b0010100000xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = `_MEM_TYPE_BYTE;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd1;
                inst_string = {8'd108 ,8'd100 ,8'd46 ,8'd98}; //ld.b
            end
            32'b0010100001xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = `_MEM_TYPE_HALF;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd1;
                inst_string = {8'd108 ,8'd100 ,8'd46 ,8'd104}; //ld.h
            end
            32'b0010100010xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd1;
                inst_string = {8'd108 ,8'd100 ,8'd46 ,8'd119}; //ld.w
            end
            32'b0010100100xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = `_MEM_TYPE_BYTE;
                decode_info.m1.mem_write = 1'd1;
                decode_info.m1.mem_valid = 1'd1;
                inst_string = {8'd115 ,8'd116 ,8'd46 ,8'd98}; //st.b
            end
            32'b0010100101xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = `_MEM_TYPE_HALF;
                decode_info.m1.mem_write = 1'd1;
                decode_info.m1.mem_valid = 1'd1;
                inst_string = {8'd115 ,8'd116 ,8'd46 ,8'd104}; //st.h
            end
            32'b0010100110xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info.m1.mem_write = 1'd1;
                decode_info.m1.mem_valid = 1'd1;
                inst_string = {8'd115 ,8'd116 ,8'd46 ,8'd119}; //st.w
            end
            32'b0010101000xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = `_MEM_TYPE_UBYTE;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd1;
                inst_string = {8'd108 ,8'd100 ,8'd46 ,8'd98 ,8'd117}; //ld.bu
            end
            32'b0010101001xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = `_MEM_TYPE_UHALF;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd1;
                inst_string = {8'd108 ,8'd100 ,8'd46 ,8'd104 ,8'd117}; //ld.hu
            end
            32'b0010101010xxxxxxxxxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = `_MEM_TYPE_UWORD;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd1;
                inst_string = {8'd108 ,8'd100 ,8'd46 ,8'd119 ,8'd117}; //ld.wu
            end
            32'b00000000000100000xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_ADD;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd97 ,8'd100 ,8'd100 ,8'd46 ,8'd119}; //add.w
            end
            32'b00000000000100010xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_SUB;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd117 ,8'd98 ,8'd46 ,8'd119}; //sub.w
            end
            32'b00000000000100100xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd108 ,8'd116}; //slt
            end
            32'b00000000000100101xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd1;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd108 ,8'd116 ,8'd117}; //sltu
            end
            32'b00000000000101000xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_NOR;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd110 ,8'd111 ,8'd114}; //nor
            end
            32'b00000000000101001xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_AND;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd97 ,8'd110 ,8'd100}; //and
            end
            32'b00000000000101010xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_OR;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd111 ,8'd114}; //or
            end
            32'b00000000000101011xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_XOR;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd120 ,8'd111 ,8'd114}; //xor
            end
            32'b00000000000101110xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_SL;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd108 ,8'd108 ,8'd46 ,8'd119}; //sll.w
            end
            32'b00000000000101111xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_SR;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd1;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd114 ,8'd108 ,8'd46 ,8'd119}; //srl.w
            end
            32'b00000000000110000xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_SR;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd114 ,8'd97 ,8'd46 ,8'd119}; //sra.w
            end
            32'b00000000000111000xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_MUL;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd109 ,8'd117 ,8'd108 ,8'd46 ,8'd119}; //mul.w
            end
            32'b00000000000111001xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_MULH;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd109 ,8'd117 ,8'd108 ,8'd104 ,8'd46 ,8'd119}; //mulh.w
            end
            32'b00000000000111010xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_MULH;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd1;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd109 ,8'd117 ,8'd108 ,8'd104 ,8'd46 ,8'd119 ,8'd117}; //mulh.wu
            end
            32'b00000000001000000xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_DIV;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd100 ,8'd105 ,8'd118 ,8'd46 ,8'd119}; //div.w
            end
            32'b00000000001000001xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_MOD;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd109 ,8'd111 ,8'd100 ,8'd46 ,8'd119}; //mod.w
            end
            32'b00000000001000010xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_DIV;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd1;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd100 ,8'd105 ,8'd118 ,8'd46 ,8'd119 ,8'd117}; //div.wu
            end
            32'b00000000001000011xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_MOD;
                decode_info.ex.opd_type = `_OPD_REG;
                decode_info.ex.opd_unsigned = 1'd1;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd109 ,8'd111 ,8'd100 ,8'd46 ,8'd119 ,8'd117}; //mod.wu
            end
            32'b00000000001010100xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RRW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd98 ,8'd114 ,8'd101 ,8'd97 ,8'd107}; //break
            end
            32'b00000000001010110xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RRW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd121 ,8'd115 ,8'd99 ,8'd97 ,8'd108 ,8'd108}; //syscall
            end
            32'b00000000010000001xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_SL;
                decode_info.ex.opd_type = `_OPD_IMM_U5;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd108 ,8'd108 ,8'd105 ,8'd46 ,8'd119}; //slli.w
            end
            32'b00000000010001001xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_SR;
                decode_info.ex.opd_type = `_OPD_IMM_U5;
                decode_info.ex.opd_unsigned = 1'd1;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd114 ,8'd108 ,8'd105 ,8'd46 ,8'd119}; //srli.w
            end
            32'b00000000010010001xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = `_ALU_TYPE_SR;
                decode_info.ex.opd_type = `_OPD_IMM_U5;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd115 ,8'd114 ,8'd97 ,8'd105 ,8'd46 ,8'd119}; //srai.w
            end
            32'b00000110010010001xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RRW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd105 ,8'd100 ,8'd108 ,8'd101}; //idle
            end
            32'b00000110010010011xxxxxxxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd1;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_M2,`_USE_M2};
                decode_info.is.reg_type = `_REG_TYPE_RRW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd105 ,8'd110 ,8'd118 ,8'd116 ,8'd108 ,8'd98}; //invtlb
            end
            32'b0000000000000000011000xxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd1;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd114 ,8'd100 ,8'd99 ,8'd110 ,8'd116 ,8'd105 ,8'd100 ,8'd46 ,8'd119}; //rdcntid.w
            end
            32'b0000000000000000011000xxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_LOW;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd114 ,8'd100 ,8'd99 ,8'd110 ,8'd116 ,8'd118 ,8'd108 ,8'd46 ,8'd119}; //rdcntvl.w
            end
            32'b0000000000000000011001xxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_HIGH;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd114 ,8'd100 ,8'd99 ,8'd110 ,8'd116 ,8'd118 ,8'd104 ,8'd46 ,8'd119}; //rdcntvh.w
            end
            32'b0000011001001000001010xxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd1;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd116 ,8'd108 ,8'd98 ,8'd115 ,8'd114 ,8'd99 ,8'd104}; //tlbsrch
            end
            32'b0000011001001000001011xxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd1;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd116 ,8'd108 ,8'd98 ,8'd114 ,8'd100}; //tlbrd
            end
            32'b0000011001001000001100xxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd1;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd116 ,8'd108 ,8'd98 ,8'd119 ,8'd114}; //tlbwr
            end
            32'b0000011001001000001101xxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd1;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd116 ,8'd108 ,8'd98 ,8'd102 ,8'd105 ,8'd108 ,8'd108}; //tlbfill
            end
            32'b0000011001001000001110xxxxxxxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd101 ,8'd114 ,8'd116 ,8'd110}; //ertn
            end
            32'b00000100xxxxxxxxxxxxxx00000xxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd1;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd0;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info.is.reg_type = `_REG_TYPE_RW;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd99 ,8'd115 ,8'd114 ,8'd114 ,8'd100}; //csrrd
            end
            32'b00000100xxxxxxxxxxxxxx00001xxxxx: begin
                decode_info.general.inst25_0 = inst[25:0];
                decode_info.ex.alu_type = 4'd0;
                decode_info.ex.opd_type = 3'd0;
                decode_info.ex.opd_unsigned = 1'd0;
                decode_info.ex.branch_type = 2'd0;
                decode_info.ex.cmp_type = 3'd0;
                decode_info.wb.rdcntv_type = `RDCNTV_TYPE_NONE;
                decode_info.wb.do_rdcntid = 1'd0;
                decode_info.wb.do_csrrd = 1'd0;
                decode_info.m2.csr_num = 14'd0;
                decode_info.m2.csr_write_en = 1'd1;
                decode_info.m2.tlbsrch_en = 1'd0;
                decode_info.m2.tlbrd_en = 1'd0;
                decode_info.m1.tlbwr_en = 1'd0;
                decode_info.m1.tlbfill_en = 1'd0;
                decode_info.m1.invtlb_en = 1'd0;
                decode_info.is.ready_time = `_READY_M2;
                decode_info.is.use_time = {`_USE_M2,`_USE_M2};
                decode_info.is.reg_type = `_REG_TYPE_RR;
                decode_info.m1.mem_type = 3'd0;
                decode_info.m1.mem_write = 1'd0;
                decode_info.m1.mem_valid = 1'd0;
                inst_string = {8'd99 ,8'd115 ,8'd114 ,8'd119 ,8'd114}; //csrwr
            end
        endcase
    end

endmodule
