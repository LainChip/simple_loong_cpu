`include "common.svh"
`include "pipeline.svh"

module cpu_core(
    input clk,
    input rst_n,
    input [7:0] int_i,
    AXI_BUS.Slave mem_bus
);

    

endmodule