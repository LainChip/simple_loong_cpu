`ifndef _CSR_HEADER
`define _CSR_HEADER

`include "common.svh"

