`include "common.svh"
`include "decoder.svh"

module decoder(
    input logic[31:0] inst_i,
    input logic fetch_err_i,
    output decode_info_t decode_info_o,
    output logic[31:0][7:0] inst_string_o
);

    always_comb begin
        unique casez(inst_i)
            32'b010011??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_BPF;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = `_USE_EX;
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = `_BRANCH_INDIRECT;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //jirl
            end
            32'b010100??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                decode_info_o.ex.branch_type = `_BRANCH_IMMEDIATE;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //b
            end
            32'b010101??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_BPF;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_BL;
                decode_info_o.ex.branch_type = `_BRANCH_IMMEDIATE;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd1;
                inst_string_o = '0; //bl
            end
            32'b010110??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_EQL;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //beq
            end
            32'b010111??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_NEQ;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //bne
            end
            32'b011000??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_LSS;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //blt
            end
            32'b011001??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_GEQ;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //bge
            end
            32'b011010??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_LTU;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //bltu
            end
            32'b011011??????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX, `_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                decode_info_o.ex.branch_type = `_BRANCH_CONDITION;
                decode_info_o.ex.cmp_type = `_CMP_GEU;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //bgeu
            end
            32'b0001010?????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_LUI;
                decode_info_o.ex.opd_type = `_OPD_IMM_S20;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_W;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //lu12i.w
            end
            32'b0001110?????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_ADD;
                decode_info_o.ex.opd_type = `_OPD_IMM_S20;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_W;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //pcaddu12i
            end
            32'b00000100????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd1;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd1;
                decode_info_o.m2.refetch = 1'd1;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_CSR;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_M2,`_USE_M2};
                decode_info_o.is.reg_type = `_REG_TYPE_CSRXCHG;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //csrwrxchg
            end
            32'b00100000????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.m2.llsc = 1'd1;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //ll.w
            end
            32'b00100001????????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info_o.m1.mem_write = 1'd1;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.m2.llsc = 1'd1;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_CSRXCHG;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //sc.w
            end
            32'b0000001000??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info_o.ex.opd_type = `_OPD_IMM_S12;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //slti
            end
            32'b0000001001??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info_o.ex.opd_type = `_OPD_IMM_S12;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //sltui
            end
            32'b0000001010??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_ADD;
                decode_info_o.ex.opd_type = `_OPD_IMM_S12;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //addi.w
            end
            32'b0000001101??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_AND;
                decode_info_o.ex.opd_type = `_OPD_IMM_U12;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //andi
            end
            32'b0000001110??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_OR;
                decode_info_o.ex.opd_type = `_OPD_IMM_U12;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //ori
            end
            32'b0000001111??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_XOR;
                decode_info_o.ex.opd_type = `_OPD_IMM_U12;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //xori
            end
            32'b0000011000??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd1;
                decode_info_o.m2.refetch = 1'd1;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_BYTE;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd1;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //cacop
            end
            32'b0010100000??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_BYTE;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //ld.b
            end
            32'b0010100001??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_HALF;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //ld.h
            end
            32'b0010100010??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //ld.w
            end
            32'b0010100100??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_BYTE;
                decode_info_o.m1.mem_write = 1'd1;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //st.b
            end
            32'b0010100101??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_HALF;
                decode_info_o.m1.mem_write = 1'd1;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //st.h
            end
            32'b0010100110??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_WORD;
                decode_info_o.m1.mem_write = 1'd1;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RR;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //st.w
            end
            32'b0010101000??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_UBYTE;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //ld.bu
            end
            32'b0010101001??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = `_MEM_TYPE_UHALF;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd1;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_LSU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //ld.hu
            end
            32'b0010101011??????????????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //preld_nop
            end
            32'b00000000000100000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_ADD;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //add.w
            end
            32'b00000000000100010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_SUB;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //sub.w
            end
            32'b00000000000100100???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //slt
            end
            32'b00000000000100101???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_SLT;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //sltu
            end
            32'b00000000000101000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_NOR;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //nor
            end
            32'b00000000000101001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_AND;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //and
            end
            32'b00000000000101010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_OR;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //or
            end
            32'b00000000000101011???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_XOR;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //xor
            end
            32'b00000000000101110???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_SL;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //sll.w
            end
            32'b00000000000101111???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_SR;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //srl.w
            end
            32'b00000000000110000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_SR;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //sra.w
            end
            32'b00000000000111000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_MUL;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = !fetch_err_i;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //mul.w
            end
            32'b00000000000111001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_MULH;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = !fetch_err_i;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //mulh.w
            end
            32'b00000000000111010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_MULH;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = !fetch_err_i;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //mulh.wu
            end
            32'b00000000001000000???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_DIV;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = !fetch_err_i;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //div.w
            end
            32'b00000000001000001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_MOD;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = !fetch_err_i;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //mod.w
            end
            32'b00000000001000010???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_DIV;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = !fetch_err_i;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //div.wu
            end
            32'b00000000001000011???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_MOD;
                decode_info_o.ex.opd_type = `_OPD_REG;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_MDU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = !fetch_err_i;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RRW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //mod.wu
            end
            32'b00000000001010100???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_SYSCALL;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //break
            end
            32'b00000000001010110???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_SYSCALL;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //syscall
            end
            32'b00000000010000001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_SL;
                decode_info_o.ex.opd_type = `_OPD_IMM_U5;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //slli.w
            end
            32'b00000000010001001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_SR;
                decode_info_o.ex.opd_type = `_OPD_IMM_U5;
                decode_info_o.ex.opd_unsigned = 1'd1;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //srli.w
            end
            32'b00000000010010001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = `_ALU_TYPE_SR;
                decode_info_o.ex.opd_type = `_OPD_IMM_U5;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = fetch_err_i;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //srai.w
            end
            32'b00000110010010001???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd1;
                decode_info_o.m2.refetch = 1'd1;
                decode_info_o.m2.wait_hint = 1'd1;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //idle
            end
            32'b00000110010010011???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd1;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd1;
                decode_info_o.m2.refetch = 1'd1;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_M2,`_USE_M2};
                decode_info_o.is.reg_type = `_REG_TYPE_INVTLB;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //invtlb
            end
            32'b00111000011100100???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd1;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //dbar
            end
            32'b00111000011100101???????????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd1;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //ibar
            end
            32'b000000000000000001100???????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_CSR;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RDCNTID;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //rdcnt.w
            end
            32'b0000011001001000001010??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd1;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd1;
                decode_info_o.m2.refetch = 1'd1;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //tlbsrch
            end
            32'b0000011001001000001011??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd1;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd1;
                decode_info_o.m2.refetch = 1'd1;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //tlbrd
            end
            32'b0000011001001000001100??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd1;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd1;
                decode_info_o.m2.refetch = 1'd1;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //tlbwr
            end
            32'b0000011001001000001101??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd1;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd1;
                decode_info_o.m2.refetch = 1'd1;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_RW;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //tlbfill
            end
            32'b0000011001001000001110??????????: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_NONE;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd1;
                decode_info_o.m2.priv_inst = 1'd1;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'd1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_M2;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = `_REG_TYPE_I;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = '0; //ertn
            end
            default: begin
                decode_info_o.general.inst25_0 = inst_i[25:0];
                decode_info_o.ex.alu_type = 4'd0;
                decode_info_o.ex.opd_type = 3'd0;
                decode_info_o.ex.opd_unsigned = 1'd0;
                decode_info_o.m2.exception_hint = `_EXCEPTION_HINT_INVALID;
                decode_info_o.m2.do_rdcntid = 1'd0;
                decode_info_o.m2.csr_num = 14'd0;
                decode_info_o.m2.csr_write_en = 1'd0;
                decode_info_o.m2.tlbsrch_en = 1'd0;
                decode_info_o.m2.tlbrd_en = 1'd0;
                decode_info_o.m2.tlbwr_en = 1'd0;
                decode_info_o.m2.tlbfill_en = 1'd0;
                decode_info_o.m2.invtlb_en = 1'd0;
                decode_info_o.m2.do_ertn = 1'd0;
                decode_info_o.m2.priv_inst = 1'd0;
                decode_info_o.m2.refetch = 1'd0;
                decode_info_o.m2.wait_hint = 1'd0;
                decode_info_o.m1.mem_type = 3'd0;
                decode_info_o.m1.mem_write = 1'd0;
                decode_info_o.m1.mem_valid = 1'd0;
                decode_info_o.m2.llsc = 1'd0;
                decode_info_o.m2.cacop = 1'd0;
                decode_info_o.wb.debug_inst = inst_i;
                decode_info_o.wb.valid = 1'b1;
                decode_info_o.wb.wb_sel = `_REG_WB_ALU;
                decode_info_o.is.pipe_one_inst = 1'b1;
                decode_info_o.is.pipe_two_inst = 1'b0;
                decode_info_o.is.ready_time = `_READY_EX;
                decode_info_o.is.use_time = {`_USE_EX,`_USE_EX};
                decode_info_o.is.reg_type = 5'b11111;
                decode_info_o.ex.branch_type = 2'd0;
                decode_info_o.ex.cmp_type = 3'd0;
                decode_info_o.ex.branch_link = 1'd0;
                inst_string_o = {8'd78 ,8'd79 ,8'd78 ,8'd69 ,8'd86 ,8'd65 ,8'd76 ,8'd73 ,8'd68}; //NONEVALID
            end
        endcase
    end

endmodule
